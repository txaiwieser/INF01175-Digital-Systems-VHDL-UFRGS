LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY mem_rom IS
	PORT(
			entrada: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
			saida: OUT STD_LOGIC_VECTOR (7 DOWNTO 0));
END mem_rom;

ARCHITECTURE circ1 OF mem_rom IS
BEGIN
	WITH entrada SELECT
	saida <=
				"00100000" WHEN "00000000",
				"10000000" WHEN "00000001",
				"10000000" WHEN "00000010",
				"00001001" WHEN "00000011",
				"00000000" WHEN "00000100",
				"00110000" WHEN "00000101",
				"10000001" WHEN "00000110",
				"10010000" WHEN "00000111",
				"00000101" WHEN "00001000",
				"01100000" WHEN "00001001",
				"01000000" WHEN "00001010",
				"10000010" WHEN "00001011",
				"01010000" WHEN "00001100",
				"10000011" WHEN "00001101",
				"00110000" WHEN "00001110",
				"10000100" WHEN "00001111",
				"10100000" WHEN "00010000",
				"00000101" WHEN "00010001",
				--"00000000" WHEN "00010011",

				"11010000" WHEN "00010010",
				"11000000" WHEN "00010011",
				"10110000" WHEN "00010100",
				"10000110" WHEN "00010101",
				"11110000" WHEN "00010110",


				"10101010" WHEN "10000000",
				"10010010" WHEN "10000001",
				"00101000" WHEN "10000010",
				"10100111" WHEN "10000011",
				"11011011" WHEN "10000100",
				"11111100" WHEN "10000101",
				"00000010" WHEN "10000110",


				"00000000" WHEN OTHERS;


END circ1;
